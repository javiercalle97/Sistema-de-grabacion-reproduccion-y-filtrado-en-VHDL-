----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 21.11.2018 11:29:21
-- Design Name: 
-- Module Name: audio_interface - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use work.DSED.all;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity audio_interface is

    Port ( clk_12megas : in STD_LOGIC;
           reset : in STD_LOGIC;
           record_enable : in STD_LOGIC;
           sample_out : out STD_LOGIC_VECTOR (sample_size-1 downto 0);
           sample_out_ready : out STD_LOGIC;
           micro_clk : out STD_LOGIC;
           micro_data : in STD_LOGIC;
           micro_LR : out STD_LOGIC;
           play_enable : in STD_LOGIC;
           sample_in : in STD_LOGIC_VECTOR (sample_size-1 downto 0);
           sample_request : out STD_LOGIC;
           jack_sd : out STD_LOGIC;
           jack_pwd : out STD_LOGIC);
end audio_interface;



architecture Behavioral of audio_interface is

signal clk_3megas, en_2_cycles, en_4_cycles, pwm_pulse, sample_out_ready_aux, control_audio, control_micro: std_logic;

signal sample_out_aux : STD_LOGIC_VECTOR (sample_size-1 downto 0);

component relojes is
    Port ( clk_12megas : in STD_LOGIC;
           reset : in STD_LOGIC;
           clk_3megas : out STD_LOGIC;
           en_2_cycles : out STD_LOGIC;
           en_4_cycles : out STD_LOGIC);
end component;

component FSMD_microphone is
  
Port ( clk_12megas : in STD_LOGIC;
       en_4_cycles : in STD_LOGIC;
       micro_data : in STD_LOGIC;
       reset : in STD_LOGIC;
       sample_out : out STD_LOGIC_VECTOR (sample_size-1 downto 0);
       sample_out_ready : out STD_LOGIC);
end component;

component pwm is
    Port ( clk_12megas : in STD_LOGIC;
           reset : in STD_LOGIC;
           en_2_cycles : in STD_LOGIC;
           sample_in : in STD_LOGIC_VECTOR (sample_size-1 downto 0);
           sample_request : out STD_LOGIC;
           pwm_pulse : out STD_LOGIC);
           
 end component;          
begin

DUT1: relojes 
    port map (clk_12megas => clk_12megas,
           reset =>reset,
           clk_3megas => clk_3megas,
           en_2_cycles => en_2_cycles,
           en_4_cycles => en_4_cycles);
           
 DUT2: FSMD_microphone 
 port map ( clk_12megas =>clk_12megas,
       en_4_cycles => control_micro,
       micro_data => micro_data,
       reset =>reset,
       sample_out => sample_out_aux,
       sample_out_ready => sample_out_ready_aux);

DUT3:  pwm 
    Port map ( clk_12megas =>clk_12megas,
           reset =>reset,
           en_2_cycles =>control_audio,
           sample_in => sample_in,
           sample_request => sample_request, 
           pwm_pulse => pwm_pulse);
           
           
    micro_clk<=clk_3megas;
    sample_out<=sample_out_aux;
    sample_out_ready<=sample_out_ready_aux;
    micro_LR<='0';
    jack_sd<='1';
  
    jack_pwd<=pwm_pulse;
    control_micro<=en_4_cycles and record_enable;
    control_audio<=en_2_cycles and play_enable;

end Behavioral;
